* tb_magic_inv.sp
*.lib ~/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.lib ~/.volare/volare/sky130/versions/933e5f2b8e42c5ec25b83c6d242455ada6f3e926/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include test_sram.spice

V_1V8	VDD 0 DC 1.8
V_0V9	VDD2 0 DC 0.9

*X0	VDD 0 O B ram_cell
*V_RD_	O_ 0	DC 0   PULSE(0 1.8 100n 0.1n 0.1n 100n 200n ) 
*V_RDB	B_ 0	DC 1.8 PULSE(0 1.8 100n 0.1n 0.1n 100n 200n ) 
*C_RD_	O_ O	10p
*C_RDB	B_ B	10p

V_Prd	Prd 0	DC 0 PULSE(0 1.8 2n 0.01n 0.01n 0.9n 10n ) 
V_Pbl	Pbl 0	DC 0 PULSE(0 1.8 1n 0.01n 0.01n 0.9n 10n ) 
CO	O 0	0.1p
CB	B 0	0.1p

.NODESET V(X0.B_)=1.8 
*V(x0.B)=0V
X0	VDD 0 O B Prd	ram_cell_access
x1	VDD2 0 O B Pbl	BTL_equalizer
x2	VDD 0 O B Prd	ampli_diff

.control
op
*print V(x0.b) V(x0.o)
print all
.endc
*.tran 0.01n 100n 
*.plot VDD O O_ B B_
