.control 
echo "fichier 2"
.endc
