.control
echo "fichier 1"
.endc
