* tb_magic_inv.sp
*.lib ~/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.lib ~/.volare/volare/sky130/versions/933e5f2b8e42c5ec25b83c6d242455ada6f3e926/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include test_sram.spice

V_1V8	VDD 0 DC 1.8
V_0V9	VDD2 0 DC 0.9

*X0	VDD 0 O B ram_cell
*V_RD_	O_ 0	DC 0   PULSE(0 1.8 100n 0.1n 0.1n 100n 200n ) 
*V_RDB	B_ 0	DC 1.8 PULSE(0 1.8 100n 0.1n 0.1n 100n 200n ) 
*C_RD_	O_ O	10p
*C_RDB	B_ B	10p

V_Prd0	Prd0 0	DC 0 PULSE(0 1.8  2n 0.01n 0.01n 0.9n 80n ) 
V_Prd1	Prd1 0	DC 0 PULSE(0 1.8 12n 0.01n 0.01n 0.9n 80n ) 
V_Prd2	Prd2 0	DC 0 PULSE(0 1.8 22n 0.01n 0.01n 0.9n 80n ) 
V_Prd3	Prd3 0	DC 0 PULSE(0 1.8 32n 0.01n 0.01n 0.9n 80n ) 
V_Prd4	Prd4 0	DC 0 PULSE(0 1.8 42n 0.01n 0.01n 0.9n 80n ) 
V_Prd5	Prd5 0	DC 0 PULSE(0 1.8 52n 0.01n 0.01n 0.9n 80n ) 
V_Prd6	Prd6 0	DC 0 PULSE(0 1.8 62n 0.01n 0.01n 0.9n 80n ) 
V_Prd7	Prd7 0	DC 0 PULSE(0 1.8 72n 0.01n 0.01n 0.9n 80n ) 
V_Pbl	Pbl  0	DC 0 PULSE(0 1.8 1n 0.01n 0.01n 0.9n 10n ) 
V_Prd	Prd  0	DC 0 PULSE(0 1.8 2n 0.01n 0.01n 0.9n 10n ) 


CO	O 0	0.1p
CB	B 0	0.1p

.NODESET V(Xb00.B_)=1.8 
.NODESET V(Xb01.O_)=1.8 
.NODESET V(Xb02.B_)=1.8 
.NODESET V(Xb03.O_)=1.8 
.NODESET V(Xb04.B_)=1.8 
.NODESET V(Xb05.O_)=1.8 
.NODESET V(Xb06.B_)=1.8 
.NODESET V(Xb07.O_)=1.8 
*V(x0.B)=0V
Xb00	VDD 0 O B Prd0	ram_cell_access
Xb01	VDD 0 O B Prd1	ram_cell_access
Xb02	VDD 0 O B Prd2	ram_cell_access
Xb03	VDD 0 O B Prd3	ram_cell_access
Xb04	VDD 0 O B Prd4	ram_cell_access
Xb05	VDD 0 O B Prd5	ram_cell_access
Xb06	VDD 0 O B Prd6	ram_cell_access
Xb07	VDD 0 O B Prd7	ram_cell_access
x1	VDD2 0 O B Pbl	BTL_equalizer
x2	VDD 0 O B Prd	ampli_diff

.control
op
*print V(x0.b) V(x0.o)
print all
.endc
*.tran 0.01n 100n 
*.plot VDD O O_ B B_
